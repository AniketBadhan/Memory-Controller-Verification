/*
Author:Aniket Badhan
*/

module mc_assert();

endmodule