/*
Author:Aniket Badhan
*/

class mc_sbd;
	 task run();
		$display("MCSBD");
	 endtask
endclass 